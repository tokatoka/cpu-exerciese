`include "Types.h"

//forwarding unit
module Forward(

    input exmemRfWrEnableIn,
    input exmemRDIn,
    input idexRSIn,
    input idexRTIn,

    input memwbRfWrEnableIn,
    input memwbRDIn,
    input memwbRSIn,
    input memwbRTIn

)

endmodule