include "Types.h"

module EXMEM(


)



endmodule